module instr_mem_file(pc, out);

input [31:0] pc;
output reg [31:0] out;

reg [31:0] i0, i1, i2, i3, i4 , i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20;
reg [31:0] k[0:1999];

initial
begin


  i0 = 32'b10001110000100010000000000000000;
	//c1
  k[0] = 32'b10001110000100010000000000000000;
  k[3] = 32'b10001110000100100000000000001001;
  k[5] = 32'b00000010001100101001100000100100;

  k[7] = 32'b10001110000100010000000000000001;
  k[9] = 32'b10001110000100100000000000001100;
  k[11]= 32'b00000010001100101010000000100100;

  k[13] = 32'b10001110000100010000000000000010;
  k[15] = 32'b10001110000100100000000000001111;
  k[17] = 32'b00000010001100101010100000100100; 

  k[19] = 32'b00000010011101001011000000100000;
  k[21] = 32'b00000010110101011011100000100000;

  k[23] = 32'b10101110000101110000000000010010;

//   //c2
  
  k[24] = 32'b10001110000100010000000000000000;
  k[26] = 32'b10001110000100100000000000001010;
  k[28] = 32'b00000010001100101001100000100100;

  k[30] = 32'b10001110000100010000000000000001;
  k[32] = 32'b10001110000100100000000000001101;
  k[34]= 32'b00000010001100101010000000100100;

  k[36] = 32'b10001110000100010000000000000010;
  k[38] = 32'b10001110000100100000000000010000;
  k[40] = 32'b00000010001100101010100000100100; 

  k[42] = 32'b00000010011101001011000000100000;
  k[44] = 32'b00000010110101011011100000100000;

  k[46] = 32'b10101110000101110000000000010011;

// 	//c3

  k[48] = 32'b10001110000100010000000000000000;
  k[50] = 32'b10001110000100100000000000001011;
  k[52] = 32'b00000010001100101001100000100100;

  k[54] = 32'b10001110000100010000000000000001;
  k[56] = 32'b10001110000100100000000000001110;
  k[58]= 32'b00000010001100101010000000100100;

  k[60] = 32'b10001110000100010000000000000010;
  k[62] = 32'b10001110000100100000000000010001;
  k[64] = 32'b00000010001100101010100000100100; 

  k[66] = 32'b00000010011101001011000000100000;
  k[68] = 32'b00000010110101011011100000100000;

  k[70] = 32'b10101110000101110000000000010100;

// 	//c4
   k[72+15] = 32'b10001110000100010000000000000011;
   k[74+15] = 32'b10001110000100100000000000001001;
   k[76+15] = 32'b00000010001100101001100000100100;

   k[78+15] = 32'b10001110000100010000000000000100;
   k[80+15] = 32'b10001110000100100000000000001100;
   k[82+15]= 32'b00000010001100101010000000100100;

   k[84+15] = 32'b10001110000100010000000000000101;
   k[86+15] = 32'b10001110000100100000000000001111;
   k[88+15] = 32'b00000010001100101010100000100100; 

   k[90+15] = 32'b00000010011101001011000000100000;
   k[92+15] = 32'b00000010110101011011100000100000;

   k[94+15] = 32'b10101110000101110000000000010101;

 //   //c5
  
   k[96+15] = 32'b10001110000100010000000000000011;
   k[98+15] = 32'b10001110000100100000000000001010;
   k[100+15] = 32'b00000010001100101001100000100100;

   k[102+15] = 32'b10001110000100010000000000000100;
   k[104+15] = 32'b10001110000100100000000000001101;
   k[106+15]= 32'b00000010001100101010000000100100;

   k[108+15] = 32'b10001110000100010000000000000101;
   k[110+15] = 32'b10001110000100100000000000010000;
   k[112+15] = 32'b00000010001100101010100000100100; 

   k[114+15] = 32'b00000010011101001011000000100000;
   k[116+15] = 32'b00000010110101011011100000100000;

   k[118+15] = 32'b10101110000101110000000000010110;

 // 	//c6

   k[120+15] = 32'b10001110000100010000000000000011;
   k[122+15] = 32'b10001110000100100000000000001011;
   k[124+15] = 32'b00000010001100101001100000100100;

   k[126+15] = 32'b10001110000100010000000000000100;
   k[128+15] = 32'b10001110000100100000000000001110;
   k[130+15]= 32'b00000010001100101010000000100100;

   k[132+15] = 32'b10001110000100010000000000000101;
   k[134+15] = 32'b10001110000100100000000000010001;
   k[136+15] = 32'b00000010001100101010100000100100; 

   k[138+15] = 32'b00000010011101001011000000100000;
   k[140+15] = 32'b00000010110101011011100000100000;

   k[142+15] = 32'b10101110000101110000000000010111;

// 	//c7
   k[172+15] = 32'b10001110000100010000000000000110;
   k[174+15] = 32'b10001110000100100000000000001001;
   k[176+15] = 32'b00000010001100101001100000100100;

   k[178+15] = 32'b10001110000100010000000000000111;
   k[180+15] = 32'b10001110000100100000000000001100;
   k[182+15]= 32'b00000010001100101010000000100100;

   k[184+15] = 32'b10001110000100010000000000001000;
   k[186+15] = 32'b10001110000100100000000000001111;
   k[188+15] = 32'b00000010001100101010100000100100; 

   k[190+15] = 32'b00000010011101001011000000100000;
   k[192+15] = 32'b00000010110101011011100000100000;

   k[194+15] = 32'b10101110000101110000000000011000;

 //   //c8
  
   k[196+15] = 32'b10001110000100010000000000000110;
   k[198+15] = 32'b10001110000100100000000000001010;
   k[1100+15] = 32'b00000010001100101001100000100100;

   k[1102+15] = 32'b10001110000100010000000000000111;
   k[1104+15] = 32'b10001110000100100000000000001101;
   k[1106+15]= 32'b00000010001100101010000000100100;

   k[1108+15] = 32'b10001110000100010000000000001000;
   k[1110+15] = 32'b10001110000100100000000000010000;
   k[1112+15] = 32'b00000010001100101010100000100100; 

   k[1114+15] = 32'b00000010011101001011000000100000;
   k[1116+15] = 32'b00000010110101011011100000100000;

   k[1118+15] = 32'b10101110000101110000000000011001;

 // 	//c9

   k[1120+15] = 32'b10001110000100010000000000000110;
   k[1122+15] = 32'b10001110000100100000000000001011;
   k[1124+15] = 32'b00000010001100101001100000100100;

   k[1126+15] = 32'b10001110000100010000000000000111;
   k[1128+15] = 32'b10001110000100100000000000001110;
   k[1130+15]= 32'b00000010001100101010000000100100;

   k[1132+15] = 32'b10001110000100010000000000001000;
   k[1134+15] = 32'b10001110000100100000000000010001;
   k[1136+15] = 32'b00000010001100101010100000100100; 

   k[1138+15] = 32'b00000010011101001011000000100000;
   k[1140+15] = 32'b00000010110101011011100000100000;

   k[1142+15] = 32'b10101110000101110000000000011010;

end

always @(pc)
begin
	case(pc)
		1: out = i0;
		// 2: out = i1;
		// 3: out = i2;
		// 4: out = i3;
		// 5: out = i4;
		// 6: out = i5;
		// 7: out = i6;
		// 8: out = i7;
		// 9: out = i8;
		// 10: out = i9;
		// 11: out = i10;
		// 12: out = i11;
		// 13: out = i12;
		// 14: out = i13;
		// 15: out = i14;
		// 16: out = i15;
		// 17: out = i16;
		// 18: out = i17;
		// 19: out = i18;
		// 20: out = i19;
		// 21: out = i20;
		default : out = k[pc];
	endcase
	// out=k[pc];
	// $display("skygfhuvifs",pc);
end

endmodule
